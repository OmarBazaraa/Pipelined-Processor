LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU IS
    GENERIC(n: INTEGER := 16);
    PORT(
        Opr     : IN  STD_LOGIC_VECTOR(  4 DOWNTO 0);

        A       : IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);
        B       : IN  STD_LOGIC_VECTOR(n-1 DOWNTO 0);

        Res1    : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);
        Res2    : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0);

        Flags   : OUT STD_LOGIC_VECTOR(  3 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE arch_ALU OF ALU IS
    
    SIGNAL FlagZ    : STD_LOGIC;
    SIGNAL FlagN    : STD_LOGIC;
    SIGNAL FlagC    : STD_LOGIC;
    SIGNAL FlagV    : STD_LOGIC;
BEGIN


END ARCHITECTURE;
